library verilog;
use verilog.vl_types.all;
entity g58_human_player_vlg_vec_tst is
end g58_human_player_vlg_vec_tst;
