library verilog;
use verilog.vl_types.all;
entity g58_play_deck_vlg_vec_tst is
end g58_play_deck_vlg_vec_tst;
