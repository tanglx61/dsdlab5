library verilog;
use verilog.vl_types.all;
entity g58_sys_ctrl_fsm_test_vlg_vec_tst is
end g58_sys_ctrl_fsm_test_vlg_vec_tst;
