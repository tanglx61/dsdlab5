library verilog;
use verilog.vl_types.all;
entity g58_comp_player_vlg_vec_tst is
end g58_comp_player_vlg_vec_tst;
