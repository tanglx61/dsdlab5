library verilog;
use verilog.vl_types.all;
entity g58_crazy8_complete_vlg_vec_tst is
end g58_crazy8_complete_vlg_vec_tst;
